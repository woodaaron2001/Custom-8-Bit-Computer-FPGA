`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    23:40:56 10/06/2022 
// Design Name: 
// Module Name:    BCDConverter 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module BCDConverter(
    input clk,
    input en,
    input [11:0] bin_d_in,
    output [15:0] bcd_d_out,
    output rdy
    );


endmodule
